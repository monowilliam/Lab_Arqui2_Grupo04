library verilog;
use verilog.vl_types.all;
entity flip_flob_lab3_vlg_vec_tst is
end flip_flob_lab3_vlg_vec_tst;

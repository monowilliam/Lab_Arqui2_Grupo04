library verilog;
use verilog.vl_types.all;
entity flip_flob_lab3_vlg_check_tst is
    port(
        Qsalida         : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end flip_flob_lab3_vlg_check_tst;
